
`include "spi_master_base.svh"
/* BASE FUNCTION and TASK
  - task     : watchdog(cycle);  // default = 1
  - task     : waitrun(cycle);   // default = 1
  - task     : init(cycle);      // default = 1
  - task     : reset(cycle);     // default = 4
  - task     : set_miso_i(value, print);
  - task     : dbg_mosi_o();
  - function : get_mosi_o(print);
  - task     : dbg_sck_o();
  - function : get_sck_o(print);
  - task     : dbg_cs_n_o();
  - function : get_cs_n_o(print);
  - task     : set_tx_byte_i(value, print);
  - task     : set_tx_byte_valid_i(value, print);
  - task     : dbg_ready_o();
  - function : get_ready_o(print);
  - task     : dbg_rx_byte_o();
  - function : get_rx_byte_o(print);
  - task     : dbg_rx_byte_valid_o();
  - function : get_rx_byte_valid_o(print);
*/
class spi_master_test #(
    parameter            SYS_FREQ = 100_000_000,
    parameter            SCK_FREQ = 25_000_000 
    ) extends spi_master_base #(
        .SYS_FREQ        (SYS_FREQ),
        .SCK_FREQ        (SCK_FREQ)
    );
    function new(virtual spi_master_io intf, string name = "spi_master");
        super.new(intf, name);
    endfunction

    // Macro function and tasks
    extern task tx_byte_control (bit [7:0] _tx_byte_i);
    extern task rx_byte_control ();

    // User define function and tasks

endclass

program automatic spi_master_program(spi_master_io io);
    // Parameter
    parameter            SYS_FREQ = 100_000_000;
    parameter            SCK_FREQ = 25_000_000 ;
    
    spi_master_test #(
        .SYS_FREQ        (SYS_FREQ),
        .SCK_FREQ        (SCK_FREQ)
        ) spi_master;
    initial begin
        spi_master = new(io);
        spi_master.printTop("spi_master test");
        spi_master.init();
        spi_master.reset();
        fork
            begin
                spi_master.watchdog(10000);
                spi_master.warn("User program not finished before watchdog timer");
            end
            begin
                //Unit byte transfer
		spi_master.tx_byte_control(8'hA5);
		while(!spi_master.get_ready_o(0)) begin
		    spi_master.waitrun(1);
		end
		spi_master.tx_byte_control(8'hCC);
		while(!spi_master.get_ready_o(0)) begin
		    spi_master.waitrun(1);
		end
            end
            spi_master.dbg_mosi_o();
            spi_master.dbg_sck_o();
            spi_master.dbg_cs_n_o();
            spi_master.dbg_ready_o();
            spi_master.dbg_rx_byte_o();
            spi_master.dbg_rx_byte_valid_o();
        join_any
        spi_master.printDiv();
    end

endprogram

// Autogenerated valid control

task spi_master_test::tx_byte_control (bit [7:0] _tx_byte_i);
    this.info("tx_byte_control requested");
    this.set_tx_byte_i(_tx_byte_i, 1);
    this.set_tx_byte_valid_i(1, 0);

    // Check condition
    #9;
    this.done("tx_byte_control granted");

    // display

    // finish
    @(intf.cb);
    this.set_tx_byte_i(0, 0);
    this.set_tx_byte_valid_i(0, 0);
endtask

task spi_master_test::rx_byte_control ();
    this.info("rx_byte_control requested");

    // Check condition
    while(!this.get_rx_byte_valid_o(0)) @(intf.cb);
    #9;
    this.done("rx_byte_control granted");

    // display
    this.get_rx_byte_o(1);

    // finish
    @(intf.cb);
endtask
